
`define BRAM_PROG_RAM 2'b00
`define BRAM_VECTOR   2'b01
`define BRAM_PROG_ROM 2'b10
